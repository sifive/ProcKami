(*
  This module defines the physical memory interface.
*)
Require Import Kami.All.
Require Import FU.
Require Import Pmp.
Require Import MemDevice.
Require Import MemTable.
Require Import List.
Import ListNotations.
Require Import BinNums.
Import BinNat.

Section pmem.
  Variable name: string.
  Variable Xlen_over_8: nat.
  Variable Rlen_over_8: nat.
  Variable mem_params : MemParamsType.
  Variable supportZifencei : bool.
  Variable ty: Kind -> Type.

  Local Notation "^ x" := (name ++ "_" ++ x)%string (at level 0).
  Local Notation Rlen := (Rlen_over_8 * 8).
  Local Notation Xlen := (Xlen_over_8 * 8).
  Local Notation Data := (Bit Rlen).
  Local Notation PAddrSz := (Xlen).
  Local Notation PAddr := (Bit PAddrSz).
  Local Notation PktWithException := (PktWithException Xlen_over_8).
  Local Notation FullException := (FullException Xlen_over_8).
  Local Notation MemWrite := (MemWrite Rlen_over_8 PAddrSz).
  Local Notation mem_devices := (@mem_devices name Xlen_over_8 Rlen_over_8 mem_params ty).
  Local Notation MemTableEntry := (@MemTableEntry name Xlen_over_8 Rlen_over_8 mem_params ty).
  Local Notation mtbl_entry_addr := (@mtbl_entry_addr name Xlen_over_8 Rlen_over_8 mem_params ty).
  Local Notation sorted_mem_table := (@sorted_mem_table name Xlen_over_8 Rlen_over_8 mem_params ty).
  Local Notation DeviceTag := (@DeviceTag name Xlen_over_8 Rlen_over_8 mem_params ty).
  Local Notation pmp_check_access := (@pmp_check_access name Xlen_over_8 ty).
  Local Notation lgMemSz := (mem_params_size mem_params).

  Record MemRegion
    := {
         mem_region_width : N;
         mem_region_device : option (Fin.t (length mem_devices))
       }.

  Local Definition mem_table_regions
    (xs : list MemTableEntry)
    :  option (N * list MemRegion)%type
    := fold_left
         (fun acc x
           => match acc with
                | None => None
                | Some (start_addr, regions)
                  => let end_addr := N.add (mtbl_entry_addr x) (mtbl_entry_width x) in
                     let device_region
                       := {|
                            mem_region_width  := mtbl_entry_width x;
                            mem_region_device := mtbl_entry_device x
                          |} in
                     match N.compare start_addr (mtbl_entry_addr x) in comparison with
                       | Datatypes.Eq
                         => Some (end_addr, regions ++ [device_region])
                       | Datatypes.Lt
                         => Some (end_addr,
                              regions ++
                              [{|
                                mem_region_width := ((mtbl_entry_addr x) - start_addr);
                                mem_region_device := None
                               |};
                               device_region])
                       | _ => None
                       end
                end)
         xs (Some (0%N, [])).

  Definition mem_regions
    := match mem_table_regions sorted_mem_table with
         | Some (_, regions) => regions
         | _ => []
         end.

  Local Definition list_sum : list N -> N := fold_right N.add 0%N.

  Local Definition option_eqb (A : Type) (H : A -> A -> bool) (x y : option A) : bool
    := match x with
         | None   => match y with | None => true    | _ => false end
         | Some n => match y with | Some m => H n m | _ => false end
         end.

  Open Scope kami_expr.
  Open Scope kami_action.

  Local Definition mem_region_match
    (region_addr : N)
    (region : MemRegion)
    (paddr : PAddr @# ty)
    :  Bool @# ty
    := ($(N.to_nat region_addr) <= paddr) &&
       (paddr < $(N.to_nat (region_addr + mem_region_width region))).

  Local Definition mem_region_apply
    (k : Kind)
    (paddr : PAddr @# ty)
    (f : MemRegion -> PAddr @# ty -> ActionT ty k)
    :  ActionT ty (Maybe k)
    := snd
         (fold_left
           (fun acc region
             => (region :: (fst acc),
                 let region_addr := list_sum (map mem_region_width (fst acc)) in
                 LETA acc_result : Maybe k <- snd acc;
                 System [
                   DispString _ "[mem_region_apply] paddr: ";
                   DispHex paddr;
                   DispString _ "\n";
                   DispString _ ("[mem_region_apply] region start: " ++ nat_hex_string (N.to_nat region_addr) ++ "\n");
                   DispString _ ("[mem_region_apply] region width: " ++ nat_hex_string (N.to_nat (mem_region_width region)) ++ "\n");
                   DispString _ ("[mem_region_apply] region end: " ++ nat_hex_string (N.to_nat (region_addr + mem_region_width region)) ++ "\n")
                 ];
                 If #acc_result @% "valid" || !(mem_region_match region_addr region paddr)
                   then
                     System [DispString _ "[mem_region_apply] did not match.\n"];
                     Ret #acc_result
                   else
                     System [DispString _ "[mem_region_apply] matched.\n"];
                     LETA result
                       :  k
                       <- f region
                            ((paddr - $(N.to_nat region_addr)) +
                             ($(N.to_nat (list_sum
                                 (map mem_region_width
                                   (filter
                                     (fun prev_region
                                       => option_eqb Fin.eqb 
                                            (mem_region_device prev_region)
                                            (mem_region_device region))
                                     (fst acc)))))));
                     Ret (Valid #result : Maybe k @# ty)
                   as result;
                 Ret #result))
           mem_regions
           ([], Ret Invalid)).

  Definition checkForAccessFault
    (access_type : VmAccessType @# ty)
    (satp_mode : Bit SatpModeWidth @# ty)
    (mode : PrivMode @# ty)
    (paddr : PAddr @# ty)
    (paddr_len : Bit 4 @# ty)
    :  ActionT ty (Maybe (Pair DeviceTag PAddr))
    := LETA pmp_result
         :  Bool
         <- pmp_check_access access_type mode paddr paddr_len; 
       LET bound_result
         :  Bool
         <- mode == $MachineMode ||
            satp_mode == $SatpModeBare ||
            satp_select
              satp_mode
              (fun vm_mode
                => $0 ==
                   (paddr >> ($(vm_mode_width vm_mode)
                              : Bit (Nat.log2_up vm_mode_max_width) @# ty)));
       LETA mresult
         :  Maybe (Maybe (Pair DeviceTag PAddr))
         <- mem_region_apply
              paddr
              (fun region device_offset
                => Ret
                     (match mem_region_device region return Maybe (Pair DeviceTag PAddr) @# ty with
                       | None => Invalid
                       | Some dtag
                         => Valid (STRUCT {
                                "fst" ::=  $(proj1_sig (to_nat dtag));
                                "snd" ::= device_offset
                              } : Pair DeviceTag PAddr @# ty)
                       end));
       System [
         DispString _ "[checkForAccessFault] pmp result: ";
         DispBinary #pmp_result;
         DispString _ "\n";
         DispString _ "[checkForAccessFault] bound result: ";
         DispBinary #bound_result;
         DispString _ "\n";
         DispString _ ("[checkForAccessFault] num memory regions: " ++ nat_decimal_string (length mem_regions) ++ "\n");
         DispString _ ("[checkForAccessFault] num memory table entries: " ++ nat_decimal_string (length sorted_mem_table) ++ "\n");
         DispString _ "[checkForAccessFault] mresult result: ";
         DispBinary #mresult;
         DispString _ "\n"
       ];
       Ret
         (utila_opt_pkt
           (#mresult @% "data" @% "data")
           (#pmp_result && #bound_result && (#mresult @% "valid") && (#mresult @% "data" @% "valid"))).

  Definition mem_region_read
    (index : Fin.t mem_device_num_reads)
    (mode : PrivMode @# ty)
    (dtag : DeviceTag @# ty)
    (daddr : PAddr @# ty)
    :  ActionT ty Data
    := mem_device_apply dtag 
         (fun device => Vector.nth (mem_device_read device mode daddr) index).

  Definition mem_region_write
    (index : Fin.t mem_device_num_writes)
    (mode : PrivMode @# ty)
    (dtag : DeviceTag @# ty)
    (daddr : PAddr @# ty)
    (data : Data @# ty)
    (mask : Array Rlen_over_8 Bool @# ty) (* TODO generalize mask size? *)
    :  ActionT ty Bool
    := mem_device_apply dtag
         (fun device
           => Vector.nth
                (mem_device_write device mode
                  (STRUCT {
                     "addr" ::= daddr;
                     "data" ::= data;
                     "mask" ::= mask
                   } : MemWrite @# ty))
                index).

  Definition pMemReadReservation (addr: PAddr @# ty)
    : ActionT ty (Array Rlen_over_8 Bool)
    := Call result: Array Rlen_over_8 Bool
                          <- ^"readMemReservation" (SignExtendTruncLsb _ addr: Bit lgMemSz);
         Ret #result.

  Definition pMemWriteReservation (addr: PAddr @# ty)
             (mask rsv: Array Rlen_over_8 Bool @# ty)
    : ActionT ty Void
    := LET writeRq: WriteRqMask lgMemSz Rlen_over_8 Bool <- STRUCT { "addr" ::= SignExtendTruncLsb lgMemSz addr ;
                                                                     "data" ::= rsv ;
                                                                     "mask" ::= mask } ;
         Call ^"writeMemReservation" (#writeRq: _);
         Retv.

  Close Scope kami_action.
  Close Scope kami_expr.

End pmem.
