module _design(
  input struct packed{ logic[31:0] inst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} exception;} fetch$_return,
  input logic[31:0] read_reg_1$_return,
  input logic[31:0] read_reg_2$_return,
  input logic[31:0] read_freg_1$_return,
  input logic[31:0] read_freg_2$_return,
  input logic[31:0] read_freg_3$_return,
  input struct packed{ logic[31:0] data; logic[1:0] reservation; struct packed{ logic valid; logic[3:0] data;} exception$;} memRead$_return,
  input struct packed{ logic valid; logic[3:0] data;} memWrite$_return,

  output logic[31:0] fetch$_argument,
  output logic[4:0] read_reg_1$_argument,
  output logic[4:0] read_reg_2$_argument,
  output logic[4:0] read_freg_1$_argument,
  output logic[4:0] read_freg_2$_argument,
  output logic[4:0] read_freg_3$_argument,
  output logic[31:0] memRead$_argument,
  output struct packed{ logic[31:0] addr; logic[31:0] data;} memWrite$_argument,
  output struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_regWrite$_argument,
  output struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_fregWrite$_argument,
  output struct packed{ logic[11:0] index; logic[31:0] data;} proc_core_csrWrite$_argument,
  output logic fetch$_enable,
  output logic read_reg_1$_enable,
  output logic read_reg_2$_enable,
  output logic read_freg_1$_enable,
  output logic read_freg_2$_enable,
  output logic read_freg_3$_enable,
  output logic memRead$_enable,
  output logic memWrite$_enable,
  output logic proc_core_regWrite$_enable,
  output logic proc_core_fregWrite$_enable,
  output logic proc_core_csrWrite$_enable,


  input CLK,
  input RESET
);
  logic[31:0] proc_core_PC;

  logic[31:0] proc_core_PC$_read;
  logic proc_core_pipeline$_guard;
  logic proc_core_pipeline$_enable;
  logic[31:0] proc_core_pipeline$1;
  struct packed{ logic[31:0] inst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} exception;} proc_core_pipeline$0$2;
  struct packed{ struct packed{ logic[31:0] pc; logic[31:0] inst;} fst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} proc_core_pipeline$1$2;
  struct packed{ struct packed{ logic[31:0] pc; logic[31:0] inst;} fst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} proc_core_pipeline$2;
  struct packed{ struct packed{ logic[31:0] pc; logic[31:0] inst;} fst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} proc_core_pipeline$0$3;
  logic[31:0] proc_core_pipeline$0$0$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$0$0$0$1$3;
  logic proc_core_pipeline$1$0$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$0$0$0$1$3;
  logic proc_core_pipeline$2$0$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$2$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$2$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[0:0] proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[0:0] proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[0:0] proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[0:0] proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[0:0] proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[0:0] proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[0:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[0:0] proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[31:0] proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[1:0] proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[15:0] proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[2:0] proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$1$0$0$0$1$3;
  logic[32:0] proc_core_pipeline$0$0$0$1$3;
  struct packed{ logic valid; logic[31:0] data;} proc_core_pipeline$0$0$1$3;
  logic[0:0] proc_core_pipeline$1$0$1$3;
  struct packed{ logic valid;} proc_core_pipeline$0$1$3;
  struct packed{ logic valid; struct packed{ logic[31:0] pc; logic[31:0] inst; logic[1:0] mode; logic compressed$;} data;} proc_core_pipeline$1$3;
  struct packed{ struct packed{ logic[31:0] pc; logic[31:0] inst; logic[1:0] mode; logic compressed$;} fst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} proc_core_pipeline$3;
  logic[31:0] proc_core_pipeline$0$0$0$4;
  logic[31:0] proc_core_pipeline$0$0$4;
  logic[31:0] proc_core_pipeline$0$1$0$4;
  logic[31:0] proc_core_pipeline$1$0$4;
  logic[31:0] proc_core_pipeline$0$2$0$4;
  logic[31:0] proc_core_pipeline$2$0$4;
  logic[31:0] proc_core_pipeline$0$3$0$4;
  logic[31:0] proc_core_pipeline$3$0$4;
  logic[31:0] proc_core_pipeline$0$4$0$4;
  logic[31:0] proc_core_pipeline$4$0$4;
  struct packed{ logic[31:0] pc; logic[31:0] reg1; logic[31:0] reg2; logic[31:0] reg3; logic[31:0] inst; logic instMisalignedException$; logic memMisalignedException$; logic accessException$; logic[1:0] mode; logic compressed$;} proc_core_pipeline$0$4;
  struct packed{ struct packed{ logic[31:0] pc; logic[31:0] reg1; logic[31:0] reg2; logic[31:0] reg3; logic[31:0] inst; logic instMisalignedException$; logic memMisalignedException$; logic accessException$; logic[1:0] mode; logic compressed$;} fst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} proc_core_pipeline$4;
  logic[0:0] proc_core_pipeline$0$0$0$5;
  struct packed{ logic valid;} proc_core_pipeline$0$0$5;
  struct packed{ logic valid;} proc_core_pipeline$0$5;
  struct packed{ struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} proc_core_pipeline$5;
  logic[84:0] proc_core_pipeline$0$0$6;
  struct packed{ logic valid; struct packed{ struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} val1; struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} val2; logic[3:0] memBitMask; logic taken$; logic aq; logic rl; struct packed{ logic valid; logic[3:0] data;} exception;} data;} proc_core_pipeline$0$6;
  struct packed{ struct packed{ struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} val1; struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} val2; logic[3:0] memBitMask; logic taken$; logic aq; logic rl; struct packed{ logic valid; logic[3:0] data;} exception;} fst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} proc_core_pipeline$6;
  struct packed{ logic writeReg$; logic[31:0] data; struct packed{ logic valid; logic[3:0] data;} exception$;} proc_core_pipeline$0$7;
  struct packed{ logic writeReg$; logic[31:0] data; struct packed{ logic valid; logic[3:0] data;} exception$;} proc_core_pipeline$1$7;
  struct packed{ logic writeReg$; logic[31:0] data; struct packed{ logic valid; logic[3:0] data;} exception$;} proc_core_pipeline$2$7;
  struct packed{ logic writeReg$; logic[31:0] data; struct packed{ logic valid; logic[3:0] data;} exception$;} proc_core_pipeline$7;
  struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} proc_core_pipeline$8;
  struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} proc_core_pipeline$9;
  logic[2:0] proc_core_pipeline$10;
  logic[2:0] proc_core_pipeline$11;
  logic[31:0] proc_core_pipeline$12;
  logic[31:0] proc_core_pipeline$13;
  struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_pipeline$14;
  struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_pipeline$15;
  struct packed{ logic[11:0] index; logic[31:0] data;} proc_core_pipeline$16;
  logic[31:0] proc_core_pipeline$proc_core_PC$_write;
  logic[31:0] proc_core_pipeline$proc_core_PC$_read;
  logic[31:0] proc_core_PC$_write;
  logic fetch$_enable;
  logic read_reg_1$_enable;
  logic read_reg_2$_enable;
  logic read_freg_1$_enable;
  logic read_freg_2$_enable;
  logic read_freg_3$_enable;
  logic proc_core_regWrite$_enable;
  logic proc_core_fregWrite$_enable;
  logic proc_core_csrWrite$_enable;
  logic[31:0] fetch$_argument;
  logic[4:0] read_reg_1$_argument;
  logic[4:0] read_reg_2$_argument;
  logic[4:0] read_freg_1$_argument;
  logic[4:0] read_freg_2$_argument;
  logic[4:0] read_freg_3$_argument;
  struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_regWrite$_argument;
  struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_fregWrite$_argument;
  struct packed{ logic[11:0] index; logic[31:0] data;} proc_core_csrWrite$_argument;
  logic fetch$_guard;
  logic read_reg_1$_guard;
  logic read_reg_2$_guard;
  logic read_freg_1$_guard;
  logic read_freg_2$_guard;
  logic read_freg_3$_guard;
  logic proc_core_regWrite$_guard;
  logic proc_core_fregWrite$_guard;
  logic proc_core_csrWrite$_guard;

  logic[4:0] _trunc$wire$285;
  logic[15:0] _trunc$wire$233;
  logic[15:0] _trunc$wire$120;
  logic[31:0] _trunc$wire$258;
  logic[15:0] _trunc$wire$128;
  logic[15:0] _trunc$wire$136;
  struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} _trunc$wire$248;
  logic[15:0] _trunc$wire$43;
  logic[15:0] _trunc$wire$82;
  logic[34:0] _trunc$wire$262;
  logic[15:0] _trunc$wire$144;
  logic[15:0] _trunc$wire$194;
  logic[11:0] _trunc$wire$290;
  logic[11:0] _trunc$wire$149;
  logic[15:0] _trunc$wire$196;
  logic[15:0] _trunc$wire$152;
  logic[10:0] _trunc$wire$66;
  logic[15:0] _trunc$wire$84;
  logic[15:0] _trunc$wire$38;
  logic[15:0] _trunc$wire$45;
  logic[15:0] _trunc$wire$90;
  logic[11:0] _trunc$wire$33;
  logic[15:0] _trunc$wire$162;
  logic[1:0] _trunc$wire$97;
  logic[15:0] _trunc$wire$146;
  logic[15:0] _trunc$wire$200;
  logic[15:0] _trunc$wire$130;
  logic[12:0] _trunc$wire$121;
  logic[15:0] _trunc$wire$198;
  logic[15:0] _trunc$wire$154;
  logic[15:0] _trunc$wire$47;
  logic[15:0] _trunc$wire$86;
  logic[9:0] _trunc$wire$65;
  logic[15:0] _trunc$wire$138;
  logic[15:0] _trunc$wire$75;
  logic[15:0] _trunc$wire$39;
  logic[15:0] _trunc$wire$218;
  logic[35:0] _trunc$wire$261;
  logic[15:0] _trunc$wire$195;
  logic[15:0] _trunc$wire$5;
  logic[15:0] _trunc$wire$50;
  struct packed{ logic[31:0] pc; logic[31:0] inst;} _trunc$wire$2;
  logic[3:0] _trunc$wire$287;
  logic[7:0] _trunc$wire$61;
  logic[1:0] _trunc$wire$180;
  logic[15:0] _trunc$wire$32;
  logic[4:0] _trunc$wire$275;
  logic[19:0] _trunc$wire$63;
  logic[1:0] _trunc$wire$123;
  logic[15:0] _trunc$wire$174;
  logic[9:0] _trunc$wire$168;
  logic[15:0] _trunc$wire$165;
  logic[35:0] _trunc$wire$253;
  logic[11:0] _trunc$wire$266;
  struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} _trunc$wire$238;
  logic[1:0] _trunc$wire$26;
  logic[1:0] _trunc$wire$48;
  logic[1:0] _trunc$wire$193;
  logic[15:0] _trunc$wire$225;
  logic[1:0] _trunc$wire$37;
  logic[0:0] _trunc$wire$236;
  logic[15:0] _trunc$wire$99;
  logic[12:0] _trunc$wire$211;
  logic[31:0] _trunc$wire$235;
  logic[11:0] _trunc$wire$95;
  logic[6:0] _trunc$wire$9;
  logic[15:0] _trunc$wire$203;
  logic[15:0] _trunc$wire$182;
  logic[5:0] _trunc$wire$274;
  logic[15:0] _trunc$wire$88;
  logic[83:0] _trunc$wire$250;
  logic[15:0] _trunc$wire$156;
  logic[15:0] _trunc$wire$49;
  logic[11:0] _trunc$wire$219;
  logic[15:0] _trunc$wire$92;
  logic[1:0] _trunc$wire$143;
  logic[15:0] _trunc$wire$164;
  logic[11:0] _trunc$wire$101;
  logic[15:0] _trunc$wire$202;
  logic[15:0] _trunc$wire$140;
  logic[15:0] _trunc$wire$51;
  logic[15:0] _trunc$wire$11;
  logic[15:0] _trunc$wire$87;
  logic[3:0] _trunc$wire$169;
  logic[15:0] _trunc$wire$148;
  logic[15:0] _trunc$wire$105;
  logic[15:0] _trunc$wire$206;
  logic[15:0] _trunc$wire$171;
  logic[11:0] _trunc$wire$167;
  logic[1:0] _trunc$wire$270;
  logic[15:0] _trunc$wire$96;
  logic[15:0] _trunc$wire$102;
  logic[15:0] _trunc$wire$208;
  logic[15:0] _trunc$wire$175;
  logic[1:0] _trunc$wire$133;
  logic[15:0] _trunc$wire$173;
  logic[12:0] _trunc$wire$161;
  logic[15:0] _trunc$wire$215;
  logic[15:0] _trunc$wire$98;
  logic[0:0] _trunc$wire$271;
  logic[15:0] _trunc$wire$53;
  logic[15:0] _trunc$wire$199;
  logic[15:0] _trunc$wire$13;
  logic[15:0] _trunc$wire$17;
  logic[15:0] _trunc$wire$56;
  logic[34:0] _trunc$wire$257;
  logic[15:0] _trunc$wire$209;
  logic[83:0] _trunc$wire$251;
  struct packed{ logic[2:0] tag; logic[31:0] data;} _trunc$wire$289;
  logic[1:0] _trunc$wire$57;
  logic[15:0] _trunc$wire$150;
  logic[4:0] _trunc$wire$214;
  struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} _trunc$wire$245;
  logic[15:0] _trunc$wire$204;
  logic[6:0] _trunc$wire$127;
  logic[15:0] _trunc$wire$71;
  logic[10:0] _trunc$wire$170;
  logic[15:0] _trunc$wire$158;
  logic[15:0] _trunc$wire$94;
  logic[4:0] _trunc$wire$221;
  struct packed{ logic valid; logic[3:0] data;} _trunc$wire$1;
  logic[3:0] _trunc$wire$187;
  logic[11:0] _trunc$wire$213;
  logic[12:0] _trunc$wire$111;
  logic[1:0] _trunc$wire$237;
  logic[15:0] _trunc$wire$54;
  logic[15:0] _trunc$wire$178;
  logic[1:0] _trunc$wire$12;
  logic[11:0] _trunc$wire$220;
  logic[84:0] _trunc$wire$249;
  logic[1:0] _trunc$wire$91;
  logic[1:0] _trunc$wire$207;
  logic[1:0] _trunc$wire$153;
  logic[15:0] _trunc$wire$59;
  logic[2:0] _trunc$wire$62;
  logic[1:0] _trunc$wire$197;
  logic[11:0] _trunc$wire$166;
  logic[1:0] _trunc$wire$22;
  struct packed{ logic[31:0] pc; logic[31:0] inst; logic[1:0] mode; logic compressed$;} _trunc$wire$240;
  logic[1:0] _trunc$wire$44;
  logic[15:0] _trunc$wire$186;
  logic[1:0] _trunc$wire$216;
  struct packed{ logic[2:0] tag; logic[31:0] data;} _trunc$wire$288;
  logic[15:0] _trunc$wire$58;
  logic[15:0] _trunc$wire$104;
  logic[35:0] _trunc$wire$260;
  logic[15:0] _trunc$wire$177;
  logic[11:0] _trunc$wire$34;
  logic[19:0] _trunc$wire$292;
  logic[15:0] _trunc$wire$217;
  logic[15:0] _trunc$wire$160;
  logic[15:0] _trunc$wire$145;
  logic[1:0] _trunc$wire$103;
  logic[1:0] _trunc$wire$81;
  logic[34:0] _trunc$wire$256;
  logic[9:0] _trunc$wire$16;
  logic[15:0] _trunc$wire$19;
  logic[15:0] _trunc$wire$83;
  logic[6:0] _trunc$wire$157;
  logic[15:0] _trunc$wire$21;
  logic[31:0] _trunc$wire$265;
  logic[18:0] _trunc$wire$67;
  logic[31:0] _trunc$wire$3;
  logic[15:0] _trunc$wire$222;
  logic[1:0] _trunc$wire$231;
  logic[15:0] _trunc$wire$179;
  logic[15:0] _trunc$wire$100;
  logic[15:0] _trunc$wire$112;
  logic[15:0] _trunc$wire$210;
  logic[15:0] _trunc$wire$68;
  logic[1:0] _trunc$wire$18;
  logic[15:0] _trunc$wire$72;
  logic[15:0] _trunc$wire$122;
  logic[1:0] _trunc$wire$201;
  logic[15:0] _trunc$wire$183;
  logic[15:0] _trunc$wire$24;
  logic[15:0] _trunc$wire$226;
  logic[15:0] _trunc$wire$93;
  logic[1:0] _trunc$wire$227;
  logic[11:0] _trunc$wire$119;
  logic[15:0] _trunc$wire$25;
  logic[15:0] _trunc$wire$23;
  logic[19:0] _trunc$wire$64;
  logic[4:0] _trunc$wire$286;
  logic[12:0] _trunc$wire$7;
  logic[15:0] _trunc$wire$106;
  logic[8:0] _trunc$wire$60;
  logic[15:0] _trunc$wire$115;
  logic[15:0] _trunc$wire$224;
  logic[1:0] _trunc$wire$184;
  logic[4:0] _trunc$wire$42;
  logic[15:0] _trunc$wire$181;
  logic[15:0] _trunc$wire$114;
  logic[15:0] _trunc$wire$70;
  logic[1:0] _trunc$wire$189;
  logic[1:0] _trunc$wire$52;
  logic[3:0] _trunc$wire$268;
  logic[37:0] _trunc$wire$282;
  logic[12:0] _trunc$wire$205;
  logic[1:0] _trunc$wire$69;
  logic[1:0] _trunc$wire$172;
  logic[6:0] _trunc$wire$137;
  struct packed{ struct packed{ logic[31:0] pc; logic[31:0] reg1; logic[31:0] reg2; logic[31:0] reg3; logic[31:0] inst; logic instMisalignedException$; logic memMisalignedException$; logic accessException$; logic[1:0] mode; logic compressed$;} fst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} _trunc$wire$246;
  logic[12:0] _trunc$wire$151;
  struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} _trunc$wire$241;
  logic[11:0] _trunc$wire$89;
  logic[34:0] _trunc$wire$255;
  logic[15:0] _trunc$wire$14;
  logic[31:0] _trunc$wire$243;
  logic[35:0] _trunc$wire$254;
  logic[1:0] _trunc$wire$73;
  logic[1:0] _trunc$wire$113;
  logic[6:0] _trunc$wire$147;
  logic[2:0] _trunc$wire$269;
  logic[36:0] _trunc$wire$283;
  logic[15:0] _trunc$wire$135;
  logic[11:0] _trunc$wire$139;
  struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} _trunc$wire$279;
  logic[4:0] _trunc$wire$35;
  logic[15:0] _trunc$wire$20;
  logic[6:0] _trunc$wire$117;
  struct packed{ struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} val1; struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} val2; logic[3:0] memBitMask; logic taken$; logic aq; logic rl; struct packed{ logic valid; logic[3:0] data;} exception;} _trunc$wire$0;
  struct packed{ logic RV32I; logic RV64I; logic Zifencei; logic Zicsr; logic RV32M; logic RV64M; logic RV32A; logic RV64A; logic RV32F; logic RV64F; logic RV32D; logic RV64D; logic RV32C; logic RV64C;} _trunc$wire$15;
  logic[6:0] _trunc$wire$273;
  logic[12:0] _trunc$wire$131;
  logic[1:0] _trunc$wire$85;
  logic[15:0] _trunc$wire$29;
  logic[15:0] _trunc$wire$116;
  logic[5:0] _trunc$wire$8;
  logic[4:0] _trunc$wire$276;
  logic[15:0] _trunc$wire$27;
  logic[32:0] _trunc$wire$234;
  logic[15:0] _trunc$wire$74;
  logic[15:0] _trunc$wire$230;
  logic[15:0] _trunc$wire$108;
  logic[15:0] _trunc$wire$188;
  logic[15:0] _trunc$wire$124;
  logic[3:0] _trunc$wire$278;
  logic[15:0] _trunc$wire$185;
  logic[15:0] _trunc$wire$132;
  logic[24:0] _trunc$wire$293;
  logic[11:0] _trunc$wire$109;
  logic[15:0] _trunc$wire$4;
  logic[15:0] _trunc$wire$76;
  logic[15:0] _trunc$wire$228;
  logic[15:0] _trunc$wire$80;
  logic[0:0] _trunc$wire$247;
  logic[15:0] _trunc$wire$46;
  logic[15:0] _trunc$wire$155;
  logic[15:0] _trunc$wire$142;
  logic[3:0] _trunc$wire$267;
  logic[11:0] _trunc$wire$212;
  struct packed{ struct packed{ logic[31:0] pc; logic[31:0] inst; logic[1:0] mode; logic compressed$;} fst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} _trunc$wire$239;
  logic[15:0] _trunc$wire$192;
  logic[15:0] _trunc$wire$79;
  logic[7:0] _trunc$wire$272;
  logic[15:0] _trunc$wire$126;
  logic[15:0] _trunc$wire$36;
  logic[4:0] _trunc$wire$284;
  logic[15:0] _trunc$wire$232;
  logic[34:0] _trunc$wire$264;
  logic[15:0] _trunc$wire$190;
  logic[15:0] _trunc$wire$134;
  logic[11:0] _trunc$wire$159;
  struct packed{ struct packed{ struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} val1; struct packed{ logic valid; struct packed{ logic[2:0] tag; logic[31:0] data;} data;} val2; logic[3:0] memBitMask; logic taken$; logic aq; logic rl; struct packed{ logic valid; logic[3:0] data;} exception;} fst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} snd;} _trunc$wire$280;
  logic[15:0] _trunc$wire$110;
  logic[15:0] _trunc$wire$78;
  logic[15:0] _trunc$wire$191;
  logic[15:0] _trunc$wire$31;
  logic[1:0] _trunc$wire$223;
  logic[15:0] _trunc$wire$118;
  logic[15:0] _trunc$wire$28;
  logic[4:0] _trunc$wire$10;
  logic[11:0] _trunc$wire$129;
  logic[34:0] _trunc$wire$263;
  logic[83:0] _trunc$wire$252;
  logic[11:0] _trunc$wire$55;
  logic[1:0] _trunc$wire$163;
  logic[11:0] _trunc$wire$41;
  logic[11:0] _trunc$wire$40;
  logic[1:0] _trunc$wire$176;
  logic[1:0] _trunc$wire$244;
  logic[47:0] _trunc$wire$259;
  logic[15:0] _trunc$wire$125;
  logic[31:0] _trunc$wire$291;
  logic[37:0] _trunc$wire$281;
  logic[6:0] _trunc$wire$107;
  logic[1:0] _trunc$wire$77;
  logic[1:0] _trunc$wire$30;
  struct packed{ logic[3:0] exception; logic[31:0] value;} _trunc$wire$242;
  logic[10:0] _trunc$wire$6;
  logic[15:0] _trunc$wire$229;
  logic[12:0] _trunc$wire$141;
  logic[4:0] _trunc$wire$277;



  assign _trunc$wire$285 = _trunc$wire$284[4:0];
  assign _trunc$wire$233 = _trunc$wire$232[15:0];
  assign _trunc$wire$120 = proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$258 = _trunc$wire$256[31:0];
  assign _trunc$wire$128 = proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$136 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$248 = proc_core_pipeline$4.snd;
  assign _trunc$wire$43 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$82 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$262 = _trunc$wire$260[34:0];
  assign _trunc$wire$144 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$194 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$290 = _trunc$wire$243[11:0];
  assign _trunc$wire$149 = _trunc$wire$148[11:0];
  assign _trunc$wire$196 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$152 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$66 = _trunc$wire$63[10:0];
  assign _trunc$wire$84 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$38 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$45 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$90 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$33 = {7'b0000000, {_trunc$wire$9[6:5], _trunc$wire$7[12:10]}};
  assign _trunc$wire$162 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$97 = _trunc$wire$96[1:0];
  assign _trunc$wire$146 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$200 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$130 = proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$121 = _trunc$wire$120[12:0];
  assign _trunc$wire$198 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$154 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$47 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$86 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$65 = _trunc$wire$63[9:0];
  assign _trunc$wire$138 = proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$75 = _trunc$wire$74[15:0];
  assign _trunc$wire$39 = _trunc$wire$38[15:0];
  assign _trunc$wire$218 = _trunc$wire$217[15:0];
  assign _trunc$wire$261 = _trunc$wire$260[35:0];
  assign _trunc$wire$195 = _trunc$wire$194[15:0];
  assign _trunc$wire$5 = _trunc$wire$4[15:0];
  assign _trunc$wire$50 = _trunc$wire$49[15:0];
  assign _trunc$wire$2 = proc_core_pipeline$0$3.fst;
  assign _trunc$wire$287 = _trunc$wire$285[3:0];
  assign _trunc$wire$61 = _trunc$wire$5[7:0];
  assign _trunc$wire$180 = _trunc$wire$179[1:0];
  assign _trunc$wire$32 = _trunc$wire$31[15:0];
  assign _trunc$wire$275 = _trunc$wire$251[4:0];
  assign _trunc$wire$63 = {9'b000000000, {_trunc$wire$7[12:12], {_trunc$wire$60[8:8], {_trunc$wire$6[10:9], {_trunc$wire$9[6:6], {_trunc$wire$61[7:7], {_trunc$wire$62[2:2], {_trunc$wire$55[11:11], _trunc$wire$8[5:3]}}}}}}}};
  assign _trunc$wire$123 = _trunc$wire$122[1:0];
  assign _trunc$wire$174 = _trunc$wire$173[15:0];
  assign _trunc$wire$168 = _trunc$wire$166[9:0];
  assign _trunc$wire$165 = _trunc$wire$164[15:0];
  assign _trunc$wire$253 = _trunc$wire$252[83:48];
  assign _trunc$wire$266 = _trunc$wire$251[11:0];
  assign _trunc$wire$238 = proc_core_pipeline$0$3.snd;
  assign _trunc$wire$26 = _trunc$wire$25[1:0];
  assign _trunc$wire$48 = _trunc$wire$47[1:0];
  assign _trunc$wire$193 = _trunc$wire$192[1:0];
  assign _trunc$wire$225 = _trunc$wire$224[15:0];
  assign _trunc$wire$37 = _trunc$wire$36[1:0];
  assign _trunc$wire$236 = proc_core_pipeline$1$0$1$3[0:0];
  assign _trunc$wire$99 = _trunc$wire$98[15:0];
  assign _trunc$wire$211 = _trunc$wire$210[12:0];
  assign _trunc$wire$235 = proc_core_pipeline$0$0$0$1$3[31:0];
  assign _trunc$wire$95 = _trunc$wire$94[11:0];
  assign _trunc$wire$9 = _trunc$wire$5[6:0];
  assign _trunc$wire$203 = _trunc$wire$202[15:0];
  assign _trunc$wire$182 = _trunc$wire$181[15:0];
  assign _trunc$wire$274 = _trunc$wire$251[5:0];
  assign _trunc$wire$88 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$250 = proc_core_pipeline$0$0$6[83:0];
  assign _trunc$wire$156 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$49 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$219 = {6'b000000, {_trunc$wire$60[8:7], _trunc$wire$7[12:9]}};
  assign _trunc$wire$92 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$143 = _trunc$wire$142[1:0];
  assign _trunc$wire$164 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$101 = _trunc$wire$100[11:0];
  assign _trunc$wire$202 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$140 = proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$51 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$11 = proc_core_pipeline$0$0$0$1$0$0$0$0$1$3[15:0];
  assign _trunc$wire$87 = _trunc$wire$86[15:0];
  assign _trunc$wire$169 = _trunc$wire$166[3:0];
  assign _trunc$wire$148 = proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$105 = _trunc$wire$104[15:0];
  assign _trunc$wire$206 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$171 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$167 = _trunc$wire$166[11:0];
  assign _trunc$wire$270 = _trunc$wire$267[1:0];
  assign _trunc$wire$96 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$102 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$208 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$175 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$133 = _trunc$wire$132[1:0];
  assign _trunc$wire$173 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$161 = _trunc$wire$160[12:0];
  assign _trunc$wire$215 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$98 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$271 = _trunc$wire$267[0:0];
  assign _trunc$wire$53 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$199 = _trunc$wire$198[15:0];
  assign _trunc$wire$13 = proc_core_pipeline$0$0$0$1$1$0$0$0$0$1$3[15:0];
  assign _trunc$wire$17 = proc_core_pipeline$0$0$0$1$0$1$0$0$0$1$3[15:0];
  assign _trunc$wire$56 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$257 = _trunc$wire$256[34:0];
  assign _trunc$wire$209 = _trunc$wire$208[15:0];
  assign _trunc$wire$251 = _trunc$wire$250[83:0];
  assign _trunc$wire$289 = proc_core_pipeline$9.data;
  assign _trunc$wire$57 = _trunc$wire$56[1:0];
  assign _trunc$wire$150 = proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$214 = _trunc$wire$212[4:0];
  assign _trunc$wire$245 = proc_core_pipeline$3.snd;
  assign _trunc$wire$204 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$127 = _trunc$wire$126[6:0];
  assign _trunc$wire$71 = _trunc$wire$70[15:0];
  assign _trunc$wire$170 = _trunc$wire$166[10:0];
  assign _trunc$wire$158 = proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$94 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$221 = _trunc$wire$219[4:0];
  assign _trunc$wire$1 = _trunc$wire$0.exception;
  assign _trunc$wire$187 = _trunc$wire$5[3:0];
  assign _trunc$wire$213 = _trunc$wire$212[11:0];
  assign _trunc$wire$111 = _trunc$wire$110[12:0];
  assign _trunc$wire$237 = _trunc$wire$3[1:0];
  assign _trunc$wire$54 = _trunc$wire$53[15:0];
  assign _trunc$wire$178 = _trunc$wire$177[15:0];
  assign _trunc$wire$12 = _trunc$wire$11[1:0];
  assign _trunc$wire$220 = _trunc$wire$219[11:0];
  assign _trunc$wire$249 = proc_core_pipeline$0$0$6[84:0];
  assign _trunc$wire$91 = _trunc$wire$90[1:0];
  assign _trunc$wire$207 = _trunc$wire$206[1:0];
  assign _trunc$wire$153 = _trunc$wire$152[1:0];
  assign _trunc$wire$59 = _trunc$wire$58[15:0];
  assign _trunc$wire$62 = _trunc$wire$5[2:0];
  assign _trunc$wire$197 = _trunc$wire$196[1:0];
  assign _trunc$wire$166 = {4'b0000, {_trunc$wire$7[12:12], {_trunc$wire$9[6:5], {_trunc$wire$62[2:2], {_trunc$wire$55[11:10], _trunc$wire$10[4:3]}}}}};
  assign _trunc$wire$22 = _trunc$wire$21[1:0];
  assign _trunc$wire$240 = proc_core_pipeline$3.fst;
  assign _trunc$wire$44 = _trunc$wire$43[1:0];
  assign _trunc$wire$186 = _trunc$wire$185[15:0];
  assign _trunc$wire$216 = _trunc$wire$215[1:0];
  assign _trunc$wire$288 = proc_core_pipeline$8.data;
  assign _trunc$wire$58 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$104 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$260 = _trunc$wire$259[47:12];
  assign _trunc$wire$177 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$34 = _trunc$wire$33[11:0];
  assign _trunc$wire$292 = _trunc$wire$243[19:0];
  assign _trunc$wire$217 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$160 = proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$145 = _trunc$wire$144[15:0];
  assign _trunc$wire$103 = _trunc$wire$102[1:0];
  assign _trunc$wire$81 = _trunc$wire$80[1:0];
  assign _trunc$wire$256 = _trunc$wire$255[34:0];
  assign _trunc$wire$16 = _trunc$wire$5[9:0];
  assign _trunc$wire$19 = proc_core_pipeline$0$0$0$1$1$0$1$0$0$0$1$3[15:0];
  assign _trunc$wire$83 = _trunc$wire$82[15:0];
  assign _trunc$wire$157 = _trunc$wire$156[6:0];
  assign _trunc$wire$21 = proc_core_pipeline$0$0$0$1$0$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$265 = _trunc$wire$263[31:0];
  assign _trunc$wire$67 = _trunc$wire$63[18:0];
  assign _trunc$wire$3 = _trunc$wire$2.inst;
  assign _trunc$wire$222 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$231 = _trunc$wire$230[1:0];
  assign _trunc$wire$179 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$100 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$112 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$210 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$68 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$18 = _trunc$wire$17[1:0];
  assign _trunc$wire$72 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$122 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$201 = _trunc$wire$200[1:0];
  assign _trunc$wire$183 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$24 = _trunc$wire$23[15:0];
  assign _trunc$wire$226 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$93 = _trunc$wire$92[15:0];
  assign _trunc$wire$227 = _trunc$wire$226[1:0];
  assign _trunc$wire$119 = _trunc$wire$118[11:0];
  assign _trunc$wire$25 = proc_core_pipeline$0$0$0$1$0$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$23 = proc_core_pipeline$0$0$0$1$1$0$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$64 = _trunc$wire$63[19:0];
  assign _trunc$wire$286 = _trunc$wire$285[4:0];
  assign _trunc$wire$7 = _trunc$wire$5[12:0];
  assign _trunc$wire$106 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$60 = _trunc$wire$5[8:0];
  assign _trunc$wire$115 = _trunc$wire$114[15:0];
  assign _trunc$wire$224 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$184 = _trunc$wire$183[1:0];
  assign _trunc$wire$42 = _trunc$wire$40[4:0];
  assign _trunc$wire$181 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$114 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$70 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$189 = _trunc$wire$188[1:0];
  assign _trunc$wire$52 = _trunc$wire$51[1:0];
  assign _trunc$wire$268 = _trunc$wire$267[3:0];
  assign _trunc$wire$282 = _trunc$wire$281[37:0];
  assign _trunc$wire$205 = _trunc$wire$204[12:0];
  assign _trunc$wire$69 = _trunc$wire$68[1:0];
  assign _trunc$wire$172 = _trunc$wire$171[1:0];
  assign _trunc$wire$137 = _trunc$wire$136[6:0];
  assign _trunc$wire$246 = {proc_core_pipeline$0$4, (((proc_core_pipeline$0$4.instMisalignedException$ | proc_core_pipeline$0$4.memMisalignedException$ | 1'b0) | proc_core_pipeline$0$4.accessException$ | 1'b0) ? {1'b0, {4'b0000, 32'b00000000000000000000000000000000}} : {1'b1, {((proc_core_pipeline$0$4.instMisalignedException$ ? 4'b0010 : 4'b0000) | (proc_core_pipeline$0$4.memMisalignedException$ ? 4'b0100 : 4'b0000) | (proc_core_pipeline$0$4.accessException$ ? 4'b0001 : 4'b0000) | 4'b0), 32'b00000000000000000000000000000000}})};
  assign _trunc$wire$151 = _trunc$wire$150[12:0];
  assign _trunc$wire$241 = proc_core_pipeline$2.snd;
  assign _trunc$wire$89 = _trunc$wire$88[11:0];
  assign _trunc$wire$255 = _trunc$wire$253[34:0];
  assign _trunc$wire$14 = _trunc$wire$13[15:0];
  assign _trunc$wire$243 = _trunc$wire$240.inst;
  assign _trunc$wire$254 = _trunc$wire$253[35:0];
  assign _trunc$wire$73 = _trunc$wire$72[1:0];
  assign _trunc$wire$113 = _trunc$wire$112[1:0];
  assign _trunc$wire$147 = _trunc$wire$146[6:0];
  assign _trunc$wire$269 = _trunc$wire$267[2:0];
  assign _trunc$wire$283 = _trunc$wire$281[36:0];
  assign _trunc$wire$135 = _trunc$wire$134[15:0];
  assign _trunc$wire$139 = _trunc$wire$138[11:0];
  assign _trunc$wire$279 = proc_core_pipeline$5.snd;
  assign _trunc$wire$35 = _trunc$wire$33[4:0];
  assign _trunc$wire$20 = _trunc$wire$19[15:0];
  assign _trunc$wire$117 = _trunc$wire$116[6:0];
  assign _trunc$wire$0 = proc_core_pipeline$6.fst;
  assign _trunc$wire$15 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
  assign _trunc$wire$273 = _trunc$wire$251[6:0];
  assign _trunc$wire$131 = _trunc$wire$130[12:0];
  assign _trunc$wire$85 = _trunc$wire$84[1:0];
  assign _trunc$wire$29 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$116 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$8 = _trunc$wire$5[5:0];
  assign _trunc$wire$276 = _trunc$wire$275[4:0];
  assign _trunc$wire$27 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$234 = proc_core_pipeline$0$0$0$1$3[32:0];
  assign _trunc$wire$74 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$230 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$108 = proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$188 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$124 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$278 = _trunc$wire$276[3:0];
  assign _trunc$wire$185 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$132 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$293 = _trunc$wire$243[24:0];
  assign _trunc$wire$109 = _trunc$wire$108[11:0];
  assign _trunc$wire$4 = _trunc$wire$3[15:0];
  assign _trunc$wire$76 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$228 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$80 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$247 = proc_core_pipeline$0$0$0$5[0:0];
  assign _trunc$wire$46 = _trunc$wire$45[15:0];
  assign _trunc$wire$155 = _trunc$wire$154[15:0];
  assign _trunc$wire$142 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$267 = _trunc$wire$266[11:8];
  assign _trunc$wire$212 = {6'b000000, {_trunc$wire$16[9:7], _trunc$wire$7[12:10]}};
  assign _trunc$wire$239 = {proc_core_pipeline$1$3.data, (proc_core_pipeline$1$3.valid ? {1'b0, {4'b0000, 32'b00000000000000000000000000000000}} : {1'b1, {4'b0010, 32'b00000000000000000000000000000000}})};
  assign _trunc$wire$192 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$79 = _trunc$wire$78[15:0];
  assign _trunc$wire$272 = _trunc$wire$251[7:0];
  assign _trunc$wire$126 = proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$36 = proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$284 = _trunc$wire$281[4:0];
  assign _trunc$wire$232 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$264 = _trunc$wire$263[34:0];
  assign _trunc$wire$190 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$134 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$159 = _trunc$wire$158[11:0];
  assign _trunc$wire$280 = {proc_core_pipeline$0$6.data, (proc_core_pipeline$0$6.valid ? {1'b0, {4'b0000, 32'b00000000000000000000000000000000}} : {1'b1, {4'b0010, 32'b00000000000000000000000000000000}})};
  assign _trunc$wire$110 = proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$78 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$191 = _trunc$wire$190[15:0];
  assign _trunc$wire$31 = proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$223 = _trunc$wire$222[1:0];
  assign _trunc$wire$118 = proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3[15:0];
  assign _trunc$wire$28 = _trunc$wire$27[15:0];
  assign _trunc$wire$10 = _trunc$wire$5[4:0];
  assign _trunc$wire$129 = _trunc$wire$128[11:0];
  assign _trunc$wire$263 = _trunc$wire$262[34:0];
  assign _trunc$wire$252 = _trunc$wire$251[83:0];
  assign _trunc$wire$55 = _trunc$wire$5[11:0];
  assign _trunc$wire$163 = _trunc$wire$162[1:0];
  assign _trunc$wire$41 = _trunc$wire$40[11:0];
  assign _trunc$wire$40 = {7'b0000000, {_trunc$wire$8[5:5], {_trunc$wire$7[12:10], _trunc$wire$9[6:6]}}};
  assign _trunc$wire$176 = _trunc$wire$175[1:0];
  assign _trunc$wire$244 = _trunc$wire$243[1:0];
  assign _trunc$wire$259 = _trunc$wire$251[47:0];
  assign _trunc$wire$125 = _trunc$wire$124[15:0];
  assign _trunc$wire$291 = _trunc$wire$243[31:0];
  assign _trunc$wire$281 = (38'b0);
  assign _trunc$wire$107 = _trunc$wire$106[6:0];
  assign _trunc$wire$77 = _trunc$wire$76[1:0];
  assign _trunc$wire$30 = _trunc$wire$29[1:0];
  assign _trunc$wire$242 = _trunc$wire$241.data;
  assign _trunc$wire$6 = _trunc$wire$5[10:0];
  assign _trunc$wire$229 = _trunc$wire$228[15:0];
  assign _trunc$wire$141 = _trunc$wire$140[12:0];
  assign _trunc$wire$277 = _trunc$wire$276[4:0];



  assign proc_core_PC$_read = proc_core_PC;
  assign proc_core_pipeline$_guard = (fetch$_guard & read_reg_1$_guard & read_reg_2$_guard & read_freg_1$_guard & read_freg_2$_guard & read_freg_3$_guard & (( ~ ( ~ _trunc$wire$1.valid)) | (( ~ proc_core_pipeline$8.valid) | ((proc_core_pipeline$10 == 3'b000) | ((proc_core_pipeline$10 == 3'b001) ? ((( ~ ( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000))) | proc_core_regWrite$_guard | 1'b0) & 1'b1) : (((proc_core_pipeline$10 == 3'b010) ? (proc_core_fregWrite$_guard & 1'b1) : ((( ~ (proc_core_pipeline$10 == 3'b011)) | proc_core_csrWrite$_guard | 1'b0) & 1'b1)) & 1'b1)) | 1'b0) | 1'b0) | (( ~ proc_core_pipeline$9.valid) | ((proc_core_pipeline$11 == 3'b000) | ((proc_core_pipeline$11 == 3'b001) ? ((( ~ ( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000))) | proc_core_regWrite$_guard | 1'b0) & 1'b1) : (((proc_core_pipeline$11 == 3'b010) ? (proc_core_fregWrite$_guard & 1'b1) : ((( ~ (proc_core_pipeline$11 == 3'b011)) | proc_core_csrWrite$_guard | 1'b0) & 1'b1)) & 1'b1)) | 1'b0) | 1'b0) | 1'b0) & 1'b1);
  assign proc_core_pipeline$_enable = proc_core_pipeline$_guard;
  assign proc_core_pipeline$1 = proc_core_pipeline$proc_core_PC$_read;
  assign proc_core_pipeline$0$2 = fetch$_return;
  assign proc_core_pipeline$1$2 = {{proc_core_pipeline$1, proc_core_pipeline$0$2.inst}, proc_core_pipeline$0$2.exception};
  assign proc_core_pipeline$2 = proc_core_pipeline$1$2;
  assign proc_core_pipeline$0$3 = proc_core_pipeline$2;
  assign proc_core_pipeline$0$0$0$0$0$1$3 = {{4'b0000, {_trunc$wire$6[10:7], {_trunc$wire$7[12:11], {_trunc$wire$8[5:5], _trunc$wire$9[6:6]}}}}, {5'b00010, {3'b000, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0010011}}}};
  assign proc_core_pipeline$0$0$0$1$0$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$0$0$0$1$3 = _trunc$wire$12[1:0];
  assign proc_core_pipeline$0$1$0$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$0$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$0$0$0$1$3 = _trunc$wire$14[15:13];
  assign proc_core_pipeline$0$1$1$0$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$0$0$0$1$3 == 3'b000);
  assign proc_core_pipeline$1$1$1$0$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$0$0$0$1$3 = (proc_core_pipeline$0$1$0$0$0$0$1$3 & proc_core_pipeline$1$1$0$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$0$0$0$1$3 = (proc_core_pipeline$0$2$0$0$0$0$1$3 | proc_core_pipeline$1$2$0$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$0$0$0$1$3 = {(proc_core_pipeline$1$0$0$0$0$1$3 & proc_core_pipeline$2$0$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$0$0$0$1$3 = {{7'b0000000, {_trunc$wire$9[6:5], _trunc$wire$7[12:10]}}, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b011, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0000111}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$0$0$0$1$3 = _trunc$wire$18[1:0];
  assign proc_core_pipeline$0$1$0$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$0$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$0$0$0$1$3 = _trunc$wire$20[15:13];
  assign proc_core_pipeline$0$1$1$0$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$0$0$0$1$3 == 3'b001);
  assign proc_core_pipeline$1$1$1$0$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$0$0$0$1$3 = _trunc$wire$15.RV32D;
  assign proc_core_pipeline$0$1$0$2$0$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$1$0$2$0$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$2$0$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$2$0$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$2$0$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$2$0$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$0$0$0$1$3 = _trunc$wire$15.RV64D;
  assign proc_core_pipeline$0$1$0$1$2$0$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$1$0$1$2$0$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$1$2$0$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$2$0$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$2$0$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$1$2$0$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$0$0$0$1$3 = {{7'b0000000, {_trunc$wire$8[5:5], {_trunc$wire$7[12:10], _trunc$wire$9[6:6]}}}, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b010, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0000011}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$0$0$0$1$3 = _trunc$wire$22[1:0];
  assign proc_core_pipeline$0$1$0$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$0$0$0$1$3 = _trunc$wire$24[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$0$0$0$1$3 == 3'b010);
  assign proc_core_pipeline$1$1$1$0$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$0$0$0$1$3 = {{7'b0000000, {_trunc$wire$8[5:5], {_trunc$wire$7[12:10], _trunc$wire$9[6:6]}}}, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b010, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0000111}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$0$0$0$1$3 = _trunc$wire$26[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$0$0$0$1$3 = _trunc$wire$28[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$0$0$0$1$3 == 3'b011);
  assign proc_core_pipeline$1$1$1$0$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32F;
  assign proc_core_pipeline$0$1$0$2$0$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$1$0$2$0$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$2$0$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$2$0$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$2$0$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$2$0$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$0$0$0$1$3 = {{7'b0000000, {_trunc$wire$9[6:5], _trunc$wire$7[12:10]}}, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b011, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0000011}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$0$0$0$1$3 = _trunc$wire$30[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$0$0$0$1$3 = _trunc$wire$32[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$0$0$0$1$3 == 3'b011);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$0$0$0$1$3 = {_trunc$wire$34[11:5], {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b011, {_trunc$wire$35[4:0], 7'b0100111}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$37[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$39[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$0$0$0$1$3 == 3'b101);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32D;
  assign proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64D;
  assign proc_core_pipeline$0$1$0$1$2$0$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$1$0$1$2$0$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$2$0$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$2$0$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$0$0$0$1$3 = {_trunc$wire$41[11:5], {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b010, {_trunc$wire$42[4:0], 7'b0100011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$44[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$46[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$0$0$0$1$3 == 3'b110);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$0$0$0$1$3 = {_trunc$wire$41[11:5], {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b010, {_trunc$wire$42[4:0], 7'b0100111}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$48[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$50[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b111);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32F;
  assign proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = {_trunc$wire$34[11:5], {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b011, {_trunc$wire$35[4:0], 7'b0100011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$52[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$54[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b111);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{6'b000000, {_trunc$wire$7[12:12], _trunc$wire$9[6:2]}}, {_trunc$wire$55[11:7], {3'b000, {_trunc$wire$55[11:7], 7'b0010011}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$57[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$59[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b000);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{_trunc$wire$64[19:19], {_trunc$wire$65[9:0], {_trunc$wire$66[10:10], _trunc$wire$67[18:11]}}}, {5'b00001, 7'b1101111}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$69[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$71[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b001);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{6'b000000, {_trunc$wire$7[12:12], _trunc$wire$9[6:2]}}, {_trunc$wire$55[11:7], {3'b000, {_trunc$wire$55[11:7], 7'b0011011}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$73[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$75[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b001);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{6'b000000, {_trunc$wire$7[12:12], _trunc$wire$9[6:2]}}, {5'b00000, {3'b000, {_trunc$wire$55[11:7], 7'b0010011}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$77[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$79[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b010);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((_trunc$wire$55[11:7] == 5'b00010) ? {{6'b000000, {_trunc$wire$7[12:12], {_trunc$wire$10[4:3], {_trunc$wire$8[5:5], {_trunc$wire$62[2:2], _trunc$wire$9[6:6]}}}}}, {5'b00010, {3'b000, {5'b00010, 7'b0010011}}}} : {{14'b00000000000000, {_trunc$wire$7[12:12], _trunc$wire$9[6:2]}}, {_trunc$wire$55[11:7], 7'b0110111}});
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$81[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$83[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b011);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {6'b000000, {{_trunc$wire$7[12:12], _trunc$wire$9[6:2]}, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b101, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0010011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$85[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$87[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$89[11:10];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {6'b010000, {{_trunc$wire$7[12:12], _trunc$wire$9[6:2]}, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b101, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0010011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$91[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$93[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$95[11:10];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{6'b000000, {_trunc$wire$7[12:12], _trunc$wire$9[6:2]}}, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b111, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0010011}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$97[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$99[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$101[11:10];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {7'b0100000, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b000, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0110011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$103[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$105[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$107[6:5];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$109[11:10];
  assign proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b11);
  assign proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$111[12:12];
  assign proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 1'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {7'b0000000, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b100, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0110011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$113[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$115[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$117[6:5];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$119[11:10];
  assign proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b11);
  assign proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$121[12:12];
  assign proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 1'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {7'b0000000, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b110, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0110011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$123[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$125[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$127[6:5];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$129[11:10];
  assign proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b11);
  assign proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$131[12:12];
  assign proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 1'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {7'b0000000, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b111, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0110011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$133[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$135[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$137[6:5];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b11);
  assign proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$139[11:10];
  assign proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b11);
  assign proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$141[12:12];
  assign proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 1'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {7'b0100000, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b000, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0111011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$143[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$145[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$147[6:5];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b00);
  assign proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$149[11:10];
  assign proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b11);
  assign proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$151[12:12];
  assign proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 1'b1);
  assign proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {7'b0000000, {(((_trunc$wire$10[4:2] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$10[4:2] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b000, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), 7'b0111011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$153[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$155[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$157[6:5];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$159[11:10];
  assign proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b11);
  assign proc_core_pipeline$0$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$161[12:12];
  assign proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 1'b1);
  assign proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{_trunc$wire$64[19:19], {_trunc$wire$65[9:0], {_trunc$wire$66[10:10], _trunc$wire$67[18:11]}}}, {5'b00000, 7'b1101111}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$163[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$165[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b101);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{_trunc$wire$167[11:11], _trunc$wire$168[9:4]}, {5'b00000, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b000, {{_trunc$wire$169[3:0], _trunc$wire$170[10:10]}, 7'b1100011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$172[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$174[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b110);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{_trunc$wire$167[11:11], _trunc$wire$168[9:4]}, {5'b00000, {(((_trunc$wire$16[9:7] == 3'b000) ? 5'b01000 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b001) ? 5'b01001 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b010) ? 5'b01010 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b011) ? 5'b01011 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b100) ? 5'b01100 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b101) ? 5'b01101 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b110) ? 5'b01110 : 5'b00000) | ((_trunc$wire$16[9:7] == 3'b111) ? 5'b01111 : 5'b00000) | 5'b0), {3'b001, {{_trunc$wire$169[3:0], _trunc$wire$170[10:10]}, 7'b1100011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$176[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b01);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$178[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b111);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {6'b000000, {{_trunc$wire$7[12:12], _trunc$wire$9[6:2]}, {_trunc$wire$55[11:7], {3'b001, {_trunc$wire$55[11:7], 7'b0010011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$180[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$182[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b000);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{6'b000000, {_trunc$wire$10[4:2], {_trunc$wire$7[12:12], _trunc$wire$9[6:5]}}}, {5'b00010, {3'b011, {_trunc$wire$55[11:7], 7'b0000111}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$184[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$186[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b001);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32D;
  assign proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64D;
  assign proc_core_pipeline$0$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{6'b000000, {_trunc$wire$187[3:2], {_trunc$wire$7[12:12], _trunc$wire$9[6:4]}}}, {5'b00010, {3'b010, {_trunc$wire$55[11:7], 7'b0000011}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$189[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$191[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b010);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{6'b000000, {_trunc$wire$187[3:2], {_trunc$wire$7[12:12], _trunc$wire$9[6:4]}}}, {5'b00010, {3'b010, {_trunc$wire$55[11:7], 7'b0000111}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$193[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$195[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b011);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32F;
  assign proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {{6'b000000, {_trunc$wire$10[4:2], {_trunc$wire$7[12:12], _trunc$wire$9[6:5]}}}, {5'b00010, {3'b011, {_trunc$wire$55[11:7], 7'b0000011}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$197[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$199[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b011);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((_trunc$wire$9[6:2] == 5'b00000) ? {12'b000000000000, {_trunc$wire$55[11:7], {3'b000, {5'b00000, 7'b1100111}}}} : {7'b0000000, {_trunc$wire$9[6:2], {5'b00000, {3'b000, {_trunc$wire$55[11:7], 7'b0110011}}}}});
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$201[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$203[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$205[12:12];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 1'b0);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((_trunc$wire$9[6:2] == 5'b00000) ? ((_trunc$wire$55[11:7] == 5'b00000) ? {12'b000000000001, {13'b0000000000000, 7'b1110011}} : {12'b000000000000, {_trunc$wire$55[11:7], {3'b000, {5'b00001, 7'b1100111}}}}) : {7'b0000000, {_trunc$wire$9[6:2], {_trunc$wire$55[11:7], {3'b000, {_trunc$wire$55[11:7], 7'b0110011}}}}});
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$207[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$209[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b100);
  assign proc_core_pipeline$0$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$211[12:12];
  assign proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 1'b1);
  assign proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {_trunc$wire$213[11:5], {_trunc$wire$9[6:2], {5'b00010, {3'b011, {_trunc$wire$214[4:0], 7'b0100111}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$216[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$218[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b101);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32D;
  assign proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64D;
  assign proc_core_pipeline$0$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {_trunc$wire$220[11:5], {_trunc$wire$9[6:2], {5'b00010, {3'b010, {_trunc$wire$221[4:0], 7'b0100011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$223[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$225[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b110);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {_trunc$wire$220[11:5], {_trunc$wire$9[6:2], {5'b00010, {3'b010, {_trunc$wire$221[4:0], 7'b0100111}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$227[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$229[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b111);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32F;
  assign proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV32C;
  assign proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {_trunc$wire$213[11:5], {_trunc$wire$9[6:2], {5'b00010, {3'b011, {_trunc$wire$214[4:0], 7'b0100011}}}}};
  assign proc_core_pipeline$0$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$231[1:0];
  assign proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 2'b10);
  assign proc_core_pipeline$0$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$4[15:0];
  assign proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$233[15:13];
  assign proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 == 3'b111);
  assign proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = _trunc$wire$15.RV64C;
  assign proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b1;
  assign proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$1$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1);
  assign proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 1'b0;
  assign proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = (proc_core_pipeline$0$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | proc_core_pipeline$1$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 1'b0);
  assign proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = {(proc_core_pipeline$1$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & proc_core_pipeline$2$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 & 1'b1), proc_core_pipeline$0$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3};
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = 33'b000000000000000000000000000000000;
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$1$0$0$0$1$3 = ((proc_core_pipeline$0$1$0$0$0$1$3.valid ? {(proc_core_pipeline$0$1$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$1$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$0$0$0$1$3 = ((proc_core_pipeline$0$0$0$0$1$3.valid ? {(proc_core_pipeline$0$0$0$0$1$3.valid ? 1'b1 : 1'b0), proc_core_pipeline$0$0$0$0$1$3.data} : 33'b000000000000000000000000000000000) | proc_core_pipeline$1$0$0$0$1$3 | 33'b0);
  assign proc_core_pipeline$0$0$1$3 = {(_trunc$wire$234[32:32] == 1'b1), _trunc$wire$235[31:0]};
  assign proc_core_pipeline$1$0$1$3 = 1'b0;
  assign proc_core_pipeline$0$1$3 = {(_trunc$wire$236[0:0] == 1'b1)};
  assign proc_core_pipeline$1$3 = {proc_core_pipeline$0$1$3.valid, {_trunc$wire$2.pc, _trunc$wire$2.inst, 2'b00, ( ~ (_trunc$wire$237[1:0] == 2'b11))}};
  assign proc_core_pipeline$3 = (_trunc$wire$238.valid ? {_trunc$wire$239.fst, proc_core_pipeline$0$3.snd} : {proc_core_pipeline$1$3.data, (proc_core_pipeline$1$3.valid ? {1'b0, {4'b0000, 32'b00000000000000000000000000000000}} : {1'b1, {4'b0010, 32'b00000000000000000000000000000000}})});
  assign proc_core_pipeline$0$0$0$4 = read_reg_1$_return;
  assign proc_core_pipeline$0$0$4 = proc_core_pipeline$0$0$0$4;
  assign proc_core_pipeline$0$1$0$4 = read_reg_2$_return;
  assign proc_core_pipeline$1$0$4 = proc_core_pipeline$0$1$0$4;
  assign proc_core_pipeline$0$2$0$4 = read_freg_1$_return;
  assign proc_core_pipeline$2$0$4 = proc_core_pipeline$0$2$0$4;
  assign proc_core_pipeline$0$3$0$4 = read_freg_2$_return;
  assign proc_core_pipeline$3$0$4 = proc_core_pipeline$0$3$0$4;
  assign proc_core_pipeline$0$4$0$4 = read_freg_3$_return;
  assign proc_core_pipeline$4$0$4 = proc_core_pipeline$0$4$0$4;
  assign proc_core_pipeline$0$4 = {_trunc$wire$240.pc, ((1'b0 ? proc_core_pipeline$0$0$4 : 32'b00000000000000000000000000000000) | (1'b0 ? proc_core_pipeline$2$0$4 : 32'b00000000000000000000000000000000) | 32'b0), ((1'b0 ? proc_core_pipeline$1$0$4 : 32'b00000000000000000000000000000000) | (1'b0 ? proc_core_pipeline$3$0$4 : 32'b00000000000000000000000000000000) | 32'b0), (1'b0 ? proc_core_pipeline$4$0$4 : 32'b00000000000000000000000000000000), _trunc$wire$240.inst, (_trunc$wire$241.valid ? (_trunc$wire$242.exception == 4'b0000) : 1'b0), (_trunc$wire$241.valid ? (_trunc$wire$242.exception == 4'b0100) : 1'b0), (_trunc$wire$241.valid ? (_trunc$wire$242.exception == 4'b0001) : 1'b0), _trunc$wire$240.mode, ( ~ (_trunc$wire$244[1:0] == 2'b11))};
  assign proc_core_pipeline$4 = (_trunc$wire$245.valid ? {_trunc$wire$246.fst, proc_core_pipeline$3.snd} : {proc_core_pipeline$0$4, (((proc_core_pipeline$0$4.instMisalignedException$ | proc_core_pipeline$0$4.memMisalignedException$ | 1'b0) | proc_core_pipeline$0$4.accessException$ | 1'b0) ? {1'b0, {4'b0000, 32'b00000000000000000000000000000000}} : {1'b1, {((proc_core_pipeline$0$4.instMisalignedException$ ? 4'b0010 : 4'b0000) | (proc_core_pipeline$0$4.memMisalignedException$ ? 4'b0100 : 4'b0000) | (proc_core_pipeline$0$4.accessException$ ? 4'b0001 : 4'b0000) | 4'b0), 32'b00000000000000000000000000000000}})});
  assign proc_core_pipeline$0$0$0$5 = 1'b0;
  assign proc_core_pipeline$0$0$5 = {(_trunc$wire$247[0:0] == 1'b1)};
  assign proc_core_pipeline$0$5 = {proc_core_pipeline$0$0$5.valid};
  assign proc_core_pipeline$5 = (_trunc$wire$248.valid ? {proc_core_pipeline$4.snd} : {(proc_core_pipeline$0$5.valid ? {1'b0, {4'b0000, 32'b00000000000000000000000000000000}} : {1'b1, {4'b0010, 32'b00000000000000000000000000000000}})});
  assign proc_core_pipeline$0$0$6 = 85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign proc_core_pipeline$0$6 = {(_trunc$wire$249[84:84] == 1'b1), {{(_trunc$wire$254[35:35] == 1'b1), {_trunc$wire$257[34:32], _trunc$wire$258[31:0]}}, {(_trunc$wire$261[35:35] == 1'b1), {_trunc$wire$264[34:32], _trunc$wire$265[31:0]}}, {(_trunc$wire$268[3:3] == 1'b1), (_trunc$wire$269[2:2] == 1'b1), (_trunc$wire$270[1:1] == 1'b1), (_trunc$wire$271[0:0] == 1'b1)}, (_trunc$wire$272[7:7] == 1'b1), (_trunc$wire$273[6:6] == 1'b1), (_trunc$wire$274[5:5] == 1'b1), {(_trunc$wire$277[4:4] == 1'b1), _trunc$wire$278[3:0]}}};
  assign proc_core_pipeline$6 = (_trunc$wire$279.valid ? {_trunc$wire$280.fst, proc_core_pipeline$5.snd} : {proc_core_pipeline$0$6.data, (proc_core_pipeline$0$6.valid ? {1'b0, {4'b0000, 32'b00000000000000000000000000000000}} : {1'b1, {4'b0010, 32'b00000000000000000000000000000000}})});
  assign proc_core_pipeline$0$7 = {(_trunc$wire$282[37:37] == 1'b1), _trunc$wire$283[36:5], {(_trunc$wire$286[4:4] == 1'b1), _trunc$wire$287[3:0]}};
  assign proc_core_pipeline$1$7 = {1'b0, 32'b00000000000000000000000000000000, {1'b0, 4'b0000}};
  assign proc_core_pipeline$2$7 = ((_trunc$wire$240.FuncUnitTag == 0) ? proc_core_pipeline$0$7 : proc_core_pipeline$1$7);
  assign proc_core_pipeline$7 = proc_core_pipeline$2$7;
  assign proc_core_pipeline$8 = _trunc$wire$0.val1;
  assign proc_core_pipeline$9 = _trunc$wire$0.val2;
  assign proc_core_pipeline$10 = _trunc$wire$288.tag;
  assign proc_core_pipeline$11 = _trunc$wire$289.tag;
  assign proc_core_pipeline$12 = _trunc$wire$288.data;
  assign proc_core_pipeline$13 = _trunc$wire$289.data;
  assign proc_core_pipeline$14 = {_trunc$wire$290[11:7], proc_core_pipeline$12};
  assign proc_core_pipeline$15 = {_trunc$wire$290[11:7], proc_core_pipeline$13};
  assign proc_core_pipeline$16 = {_trunc$wire$291[31:20], proc_core_pipeline$13};
  assign proc_core_pipeline$proc_core_PC$_write = proc_core_pipeline$proc_core_PC$_read;
  assign proc_core_pipeline$proc_core_PC$_read = proc_core_PC$_read;
  assign proc_core_PC$_write = proc_core_pipeline$proc_core_PC$_write;
  assign fetch$_enable = (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1);
  assign read_reg_1$_enable = (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1);
  assign read_reg_2$_enable = (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1);
  assign read_freg_1$_enable = (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1);
  assign read_freg_2$_enable = (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1);
  assign read_freg_3$_enable = (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1);
  assign proc_core_regWrite$_enable = (( ~ _trunc$wire$1.valid) ? ((proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0) : 1'b0)) : 1'b0) ? (proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0) : 1'b0)) : 1'b0) : (proc_core_pipeline$8.valid ? ((proc_core_pipeline$10 == 3'b000) ? 1'b0 : ((proc_core_pipeline$10 == 3'b001) ? (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0) : 1'b0)) : 1'b0)) : 1'b0);
  assign proc_core_fregWrite$_enable = (( ~ _trunc$wire$1.valid) ? ((proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? 1'b0 : ((proc_core_pipeline$11 == 3'b010) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0))) : 1'b0) ? (proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? 1'b0 : ((proc_core_pipeline$11 == 3'b010) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0))) : 1'b0) : (proc_core_pipeline$8.valid ? ((proc_core_pipeline$10 == 3'b000) ? 1'b0 : ((proc_core_pipeline$10 == 3'b001) ? 1'b0 : ((proc_core_pipeline$10 == 3'b010) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0))) : 1'b0)) : 1'b0);
  assign proc_core_csrWrite$_enable = (( ~ _trunc$wire$1.valid) ? ((proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? 1'b0 : ((proc_core_pipeline$11 == 3'b010) ? 1'b0 : ((proc_core_pipeline$11 == 3'b011) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0)))) : 1'b0) ? (proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? 1'b0 : ((proc_core_pipeline$11 == 3'b010) ? 1'b0 : ((proc_core_pipeline$11 == 3'b011) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0)))) : 1'b0) : (proc_core_pipeline$8.valid ? ((proc_core_pipeline$10 == 3'b000) ? 1'b0 : ((proc_core_pipeline$10 == 3'b001) ? 1'b0 : ((proc_core_pipeline$10 == 3'b010) ? 1'b0 : ((proc_core_pipeline$10 == 3'b011) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0)))) : 1'b0)) : 1'b0);
  assign fetch$_argument = proc_core_pipeline$1;
  assign read_reg_1$_argument = _trunc$wire$292[19:15];
  assign read_reg_2$_argument = _trunc$wire$293[24:20];
  assign read_freg_1$_argument = _trunc$wire$292[19:15];
  assign read_freg_2$_argument = _trunc$wire$293[24:20];
  assign read_freg_3$_argument = _trunc$wire$291[31:27];
  assign proc_core_regWrite$_argument = (( ~ _trunc$wire$1.valid) ? ((proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0) : 1'b0)) : 1'b0) ? (proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15) : (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15)) : ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15) : (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15))) : ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15) : (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15)) : ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15) : (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15)))) : (proc_core_pipeline$8.valid ? ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14) : (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14)) : ((proc_core_pipeline$10 == 3'b001) ? (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14) : (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14))) : ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14) : (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14)) : ((proc_core_pipeline$10 == 3'b001) ? (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14) : (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14))))) : ((proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0) : 1'b0)) : 1'b0) ? (proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15) : (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15)) : ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15) : (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15))) : ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15) : (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15)) : ((proc_core_pipeline$11 == 3'b001) ? (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15) : (( ~ (proc_core_pipeline$15.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$15 : proc_core_pipeline$15)))) : (proc_core_pipeline$8.valid ? ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14) : (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14)) : ((proc_core_pipeline$10 == 3'b001) ? (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14) : (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14))) : ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14) : (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14)) : ((proc_core_pipeline$10 == 3'b001) ? (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14) : (( ~ (proc_core_pipeline$14.data == 32'b00000000000000000000000000000000)) ? proc_core_pipeline$14 : proc_core_pipeline$14))))));
  assign proc_core_fregWrite$_argument = (( ~ _trunc$wire$1.valid) ? ((proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? 1'b0 : ((proc_core_pipeline$11 == 3'b010) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0))) : 1'b0) ? (proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15) : ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15)) : ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15) : ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15))) : ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15) : ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15)) : ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15) : ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15)))) : (proc_core_pipeline$8.valid ? ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14) : ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14)) : ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14) : ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14))) : ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14) : ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14)) : ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14) : ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14))))) : ((proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? 1'b0 : ((proc_core_pipeline$11 == 3'b010) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0))) : 1'b0) ? (proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15) : ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15)) : ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15) : ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15))) : ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15) : ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15)) : ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15) : ((proc_core_pipeline$11 == 3'b010) ? proc_core_pipeline$15 : proc_core_pipeline$15)))) : (proc_core_pipeline$8.valid ? ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14) : ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14)) : ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14) : ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14))) : ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14) : ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14)) : ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14) : ((proc_core_pipeline$10 == 3'b010) ? proc_core_pipeline$14 : proc_core_pipeline$14))))));
  assign proc_core_csrWrite$_argument = (( ~ _trunc$wire$1.valid) ? ((proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? 1'b0 : ((proc_core_pipeline$11 == 3'b010) ? 1'b0 : ((proc_core_pipeline$11 == 3'b011) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0)))) : 1'b0) ? (proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))) : ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)))) : ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))) : ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))))) : (proc_core_pipeline$8.valid ? ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))) : ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)))) : ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))) : ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)))))) : ((proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? 1'b0 : ((proc_core_pipeline$11 == 3'b001) ? 1'b0 : ((proc_core_pipeline$11 == 3'b010) ? 1'b0 : ((proc_core_pipeline$11 == 3'b011) ? (proc_core_pipeline$_guard & proc_core_pipeline$_enable & 1'b1) : 1'b0)))) : 1'b0) ? (proc_core_pipeline$9.valid ? ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))) : ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)))) : ((proc_core_pipeline$11 == 3'b000) ? ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))) : ((proc_core_pipeline$11 == 3'b001) ? ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$11 == 3'b010) ? ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$11 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))))) : (proc_core_pipeline$8.valid ? ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))) : ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)))) : ((proc_core_pipeline$10 == 3'b000) ? ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16))) : ((proc_core_pipeline$10 == 3'b001) ? ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)) : ((proc_core_pipeline$10 == 3'b010) ? ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16) : ((proc_core_pipeline$10 == 3'b011) ? proc_core_pipeline$16 : proc_core_pipeline$16)))))));
  assign fetch$_guard = 1'b1;
  assign read_reg_1$_guard = 1'b1;
  assign read_reg_2$_guard = 1'b1;
  assign read_freg_1$_guard = 1'b1;
  assign read_freg_2$_guard = 1'b1;
  assign read_freg_3$_guard = 1'b1;
  assign proc_core_regWrite$_guard = 1'b1;
  assign proc_core_fregWrite$_guard = 1'b1;
  assign proc_core_csrWrite$_guard = 1'b1;

  always @(posedge CLK) begin
    if(RESET) begin
      proc_core_PC <= 32'b00000000000000000000000000000000;
    end
    else begin
      proc_core_PC <= proc_core_PC$_write;
    end
  end
endmodule

module top(
  input struct packed{ logic[31:0] inst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} exception;} fetch$_return,
  input logic[31:0] read_reg_1$_return,
  input logic[31:0] read_reg_2$_return,
  input logic[31:0] read_freg_1$_return,
  input logic[31:0] read_freg_2$_return,
  input logic[31:0] read_freg_3$_return,

  output logic[31:0] fetch$_argument,
  output logic[4:0] read_reg_1$_argument,
  output logic[4:0] read_reg_2$_argument,
  output logic[4:0] read_freg_1$_argument,
  output logic[4:0] read_freg_2$_argument,
  output logic[4:0] read_freg_3$_argument,
  output struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_regWrite$_argument,
  output struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_fregWrite$_argument,
  output struct packed{ logic[11:0] index; logic[31:0] data;} proc_core_csrWrite$_argument,
  output logic fetch$_enable,
  output logic read_reg_1$_enable,
  output logic read_reg_2$_enable,
  output logic read_freg_1$_enable,
  output logic read_freg_2$_enable,
  output logic read_freg_3$_enable,
  output logic proc_core_regWrite$_enable,
  output logic proc_core_fregWrite$_enable,
  output logic proc_core_csrWrite$_enable,
  output logic proc_core_regWrite$_enable,
  output logic proc_core_fregWrite$_enable,
  output logic proc_core_csrWrite$_enable,

  input CLK,
  input RESET
);
  struct packed{ logic[31:0] inst; struct packed{ logic valid; struct packed{ logic[3:0] exception; logic[31:0] value;} data;} exception;} fetch$_return;
  logic[31:0] read_reg_1$_return;
  logic[31:0] read_reg_2$_return;
  logic[31:0] read_freg_1$_return;
  logic[31:0] read_freg_2$_return;
  logic[31:0] read_freg_3$_return;

  logic[31:0] fetch$_argument;
  logic[4:0] read_reg_1$_argument;
  logic[4:0] read_reg_2$_argument;
  logic[4:0] read_freg_1$_argument;
  logic[4:0] read_freg_2$_argument;
  logic[4:0] read_freg_3$_argument;
  struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_regWrite$_argument;
  struct packed{ logic[4:0] index; logic[31:0] data;} proc_core_fregWrite$_argument;
  struct packed{ logic[11:0] index; logic[31:0] data;} proc_core_csrWrite$_argument;
  logic fetch$_enable;
  logic read_reg_1$_enable;
  logic read_reg_2$_enable;
  logic read_freg_1$_enable;
  logic read_freg_2$_enable;
  logic read_freg_3$_enable;
  logic proc_core_regWrite$_enable;
  logic proc_core_fregWrite$_enable;
  logic proc_core_csrWrite$_enable;


  _design _designInst(.CLK(CLK), .RESET(RESET), .fetch$_return(fetch$_return), .read_reg_1$_return(read_reg_1$_return), .read_reg_2$_return(read_reg_2$_return), .read_freg_1$_return(read_freg_1$_return), .read_freg_2$_return(read_freg_2$_return), .read_freg_3$_return(read_freg_3$_return), .fetch$_argument(fetch$_argument), .read_reg_1$_argument(read_reg_1$_argument), .read_reg_2$_argument(read_reg_2$_argument), .read_freg_1$_argument(read_freg_1$_argument), .read_freg_2$_argument(read_freg_2$_argument), .read_freg_3$_argument(read_freg_3$_argument), .proc_core_regWrite$_argument(proc_core_regWrite$_argument), .proc_core_fregWrite$_argument(proc_core_fregWrite$_argument), .proc_core_csrWrite$_argument(proc_core_csrWrite$_argument), .fetch$_enable(fetch$_enable), .read_reg_1$_enable(read_reg_1$_enable), .read_reg_2$_enable(read_reg_2$_enable), .read_freg_1$_enable(read_freg_1$_enable), .read_freg_2$_enable(read_freg_2$_enable), .read_freg_3$_enable(read_freg_3$_enable), .proc_core_regWrite$_enable(proc_core_regWrite$_enable), .proc_core_fregWrite$_enable(proc_core_fregWrite$_enable), .proc_core_csrWrite$_enable(proc_core_csrWrite$_enable));
endmodule

